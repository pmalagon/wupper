-- ***************************************************************************
-- ***************************************************************************
-- ***************************************************************************
-- ***************************************************************************
-- ***************************************************************************
-- DO NOT EDIT THIS FILE
-- 
-- This file was generated from template '../firmware/sources/templates/register_map_sync.vhd.template'
-- and register map registers-1.0.yaml, version 2.0
-- by the script 'wuppercodegen', version: 0.8.4,
-- using the following commandline:
-- 
-- ../software/wuppercodegen/wuppercodegen/cli.py registers-1.0.yaml ../firmware/sources/templates/register_map_sync.vhd.template ../firmware/sources/pcie/register_map_sync.vhd
-- 
-- Please do NOT edit this file, but edit the source file at '../firmware/sources/templates/register_map_sync.vhd.template'
-- 
-- ***************************************************************************
-- ***************************************************************************
-- ***************************************************************************
-- ***************************************************************************
-- ***************************************************************************


--!------------------------------------------------------------------------------
--!
--!           NIKHEF - National Institute for Subatomic Physics
--!
--!                       Electronics Department
--!
--!-----------------------------------------------------------------------------
--! @class register_map_sync
--!
--!
--! @author      Andrea Borga    (andrea.borga@nikhef.nl)<br>
--!              Frans Schreuder (frans.schreuder@nikhef.nl)
--!
--!
--! @date        07/01/2015    created
--!
--! @version     1.0
--!
--! @brief
--! synchronizes the register map record to the given sync_clock
--!
--! @detail
--!
--!-----------------------------------------------------------------------------
--! @TODO
--!
--!
--! ------------------------------------------------------------------------------
--! Wupper: PCIe Gen3 and Gen4 DMA Core for Xilinx FPGAs
--! 
--! Copyright (C) 2021 Nikhef, Amsterdam (f.schreuder@nikhef.nl)
--! 
--! Licensed under the Apache License, Version 2.0 (the "License");
--! you may not use this file except in compliance with the License.
--! You may obtain a copy of the License at
--! 
--!         http://www.apache.org/licenses/LICENSE-2.0
--! 
--! Unless required by applicable law or agreed to in writing, software
--! distributed under the License is distributed on an "AS IS" BASIS,
--! WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
--! See the License for the specific language governing permissions and
--! limitations under the License.
-- 
--! @brief ieee



library ieee, UNISIM;
use ieee.numeric_std.all;
use UNISIM.VCOMPONENTS.all;
--use ieee.std_logic_unsigned.all;
use ieee.std_logic_1164.all;
use work.pcie_package.all;

entity register_map_sync is
  generic(
    NUMBER_OF_INTERRUPTS : integer := 8);
  port (
    appreg_clk                  : in     std_logic;
    clk40                       : in     std_logic;
    interrupt_call              : out    std_logic_vector(NUMBER_OF_INTERRUPTS-1 downto 4);
    interrupt_call_cr           : in     std_logic_vector(NUMBER_OF_INTERRUPTS-1 downto 4);
    register_map_40_control     : out    register_map_control_type;
    register_map_control        : in     register_map_control_type;
   register_map_gen_board_info      : in     register_map_gen_board_info_type;
   register_map_hk_monitor      : in     register_map_hk_monitor_type;
   wishbone_monitor      : in     wishbone_monitor_type;
    register_map_monitor        : out    register_map_monitor_type;
    rst_hw                      : in     std_logic;
    rst_soft_40                 : out    std_logic;
    rst_soft_appregclk          : in     std_logic;
    master_busy_in              : in     std_logic);
end entity register_map_sync;



architecture rtl of register_map_sync is

  --attribute ASYNC_REG     : string;

  --synchronization stages to 41.667MHz
  signal interrupt_call_p1                         : std_logic_vector(NUMBER_OF_INTERRUPTS-1 downto 4);

   signal register_map_gen_board_info_p1               : register_map_gen_board_info_type;
   --attribute ASYNC_REG of register_map_gen_board_info_p1            : signal is "TRUE";
   signal register_map_hk_monitor_p1               : register_map_hk_monitor_type;
   --attribute ASYNC_REG of register_map_hk_monitor_p1            : signal is "TRUE";
   signal wishbone_monitor_p1               : wishbone_monitor_type;
   --attribute ASYNC_REG of wishbone_monitor_p1            : signal is "TRUE";
  
  signal register_map_control_p1                   : register_map_control_type;
  signal rst_soft_p1                  : std_logic;
  
begin

    clk40_sync: process(clk40)
    begin
      if(rising_edge(clk40)) then
        register_map_40_control <= register_map_control_p1;
        register_map_control_p1 <= register_map_control;
        rst_soft_40 <= rst_soft_p1 or rst_hw;
        rst_soft_p1 <= rst_soft_appregclk;
      end if;
    end process;

    appreg_sync: process(appreg_clk)
      variable master_busy_p1, master_busy_p2: std_logic;
    begin
      if(rising_edge(appreg_clk)) then
        if master_busy_p1 /= master_busy_p2 then
            interrupt_call(6) <= '1';
        else 
            interrupt_call(6) <= '0';
        end if;
        
        master_busy_p2 := master_busy_p1;
        master_busy_p1 := master_busy_in;
        
      
        interrupt_call(7) <= interrupt_call_p1(7);
        interrupt_call(5) <= interrupt_call_p1(5);
        interrupt_call(4) <= interrupt_call_p1(4);
        interrupt_call_p1 <= interrupt_call_cr;
        
        register_map_monitor.register_map_gen_board_info       <= register_map_gen_board_info_p1;
        register_map_gen_board_info_p1                         <= register_map_gen_board_info;
        register_map_monitor.register_map_hk_monitor       <= register_map_hk_monitor_p1;
        register_map_hk_monitor_p1                         <= register_map_hk_monitor;
        register_map_monitor.wishbone_monitor       <= wishbone_monitor_p1;
        wishbone_monitor_p1                         <= wishbone_monitor;
        
      end if;
    end process;

end architecture rtl ; -- of register_map_sync
